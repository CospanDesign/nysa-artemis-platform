
module artemis_ddr3_user (
  input           ddr3_in_clk,
  input           rst,

  output          calibration_done,

  output          usr_clk,
  output          usr_rst,

  inout   [7:0]   mcb3_dram_dq,
  output  [13:0]  mcb3_dram_a,
  output  [2:0]   mcb3_dram_ba,
  output          mcb3_dram_ras_n,
  output          mcb3_dram_cas_n,
  output          mcb3_dram_we_n,
  output          mcb3_dram_odt,
  output          mcb3_dram_reset_n,
  output          mcb3_dram_cke,
  output          mcb3_dram_dm,
  inout           mcb3_rzq,
  inout           mcb3_zio,
  inout           mcb3_dram_dqs,
  inout           mcb3_dram_dqs_n,
  output          mcb3_dram_ck,
  output          mcb3_dram_ck_n,

  input           p0_cmd_clk,
  input           p0_cmd_en,
  input   [2:0]   p0_cmd_instr,
  input   [5:0]   p0_cmd_bl,
  input   [29:0]  p0_cmd_byte_addr,
  output          p0_cmd_empty,
  output          p0_cmd_full,
  input           p0_wr_clk,
  input           p0_wr_en,
  input   [3:0]   p0_wr_mask,
  input   [31:0]  p0_wr_data,
  output          p0_wr_full,
  output          p0_wr_empty,
  output  [6:0]   p0_wr_count,
  output          p0_wr_underrun,
  output          p0_wr_error,
  input           p0_rd_clk,
  input           p0_rd_en,
  output  [31:0]  p0_rd_data,
  output          p0_rd_full,
  output          p0_rd_empty,
  output  [6:0]   p0_rd_count,
  output          p0_rd_overflow,
  output          p0_rd_error,

  input           p1_cmd_clk,
  input           p1_cmd_en,
  input   [2:0]   p1_cmd_instr,
  input   [5:0]   p1_cmd_bl,
  input   [29:0]  p1_cmd_byte_addr,
  output          p1_cmd_empty,
  output          p1_cmd_full,
  input           p1_wr_clk,
  input           p1_wr_en,
  input   [3:0]   p1_wr_mask,
  input   [31:0]  p1_wr_data,
  output          p1_wr_full,
  output          p1_wr_empty,
  output  [6:0]   p1_wr_count,
  output          p1_wr_underrun,
  output          p1_wr_error,
  input           p1_rd_clk,
  input           p1_rd_en,
  output  [31:0]  p1_rd_data,
  output          p1_rd_full,
  output          p1_rd_empty,
  output  [6:0]   p1_rd_count,
  output          p1_rd_overflow,
  output          p1_rd_error,

  input           p2_cmd_clk,
  input           p2_cmd_en,
  input   [2:0]   p2_cmd_instr,
  input   [5:0]   p2_cmd_bl,
  input   [29:0]  p2_cmd_byte_addr,
  output          p2_cmd_empty,
  output          p2_cmd_full,
  input           p2_wr_clk,
  input           p2_wr_en,
  input   [3:0]   p2_wr_mask,
  input   [31:0]  p2_wr_data,
  output          p2_wr_full,
  output          p2_wr_empty,
  output  [6:0]   p2_wr_count,
  output          p2_wr_underrun,
  output          p2_wr_error,
  input           p2_rd_clk,
  input           p2_rd_en,
  output  [31:0]  p2_rd_data,
  output          p2_rd_full,
  output          p2_rd_empty,
  output  [6:0]   p2_rd_count,
  output          p2_rd_overflow,
  output          p2_rd_error,

  input           p3_cmd_clk,
  input           p3_cmd_en,
  input   [2:0]   p3_cmd_instr,
  input   [5:0]   p3_cmd_bl,
  input   [29:0]  p3_cmd_byte_addr,
  output          p3_cmd_empty,
  output          p3_cmd_full,
  input           p3_wr_clk,
  input           p3_wr_en,
  input   [3:0]   p3_wr_mask,
  input   [31:0]  p3_wr_data,
  output          p3_wr_full,
  output          p3_wr_empty,
  output  [6:0]   p3_wr_count,
  output          p3_wr_underrun,
  output          p3_wr_error,
  input           p3_rd_clk,
  input           p3_rd_en,
  output  [31:0]  p3_rd_data,
  output          p3_rd_full,
  output          p3_rd_empty,
  output  [6:0]   p3_rd_count,
  output          p3_rd_overflow,
  output          p3_rd_error


);
endmodule
