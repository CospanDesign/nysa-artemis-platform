

module artemis_ddr3 (
  input           clk_333mhz,
  input           board_rst,
  output          calibration_done,
  output          usr_clk,
  output          rst,

  //Memory Interface
  inout  [7:0]    ddr3_dram_dq,
  output [13:0]   ddr3_dram_a,
  output [2:0]    ddr3_dram_ba,
  output          ddr3_dram_ras_n,
  output          ddr3_dram_cas_n,
  output          ddr3_dram_we_n,
  output          ddr3_dram_odt,
  output          ddr3_dram_reset_n,
  output          ddr3_dram_cke,
  output          ddr3_dram_dm,
  inout           ddr3_rzq,
  inout           ddr3_zio,
  inout           ddr3_dram_dqs,
  inout           ddr3_dram_dqs_n,
  output          ddr3_dram_ck,
  output          ddr3_dram_ck_n,

  //Port Interfaces
  input           p0_cmd_clk,
  input           p0_cmd_en,
  input   [2:0]   p0_cmd_instr,
  input   [5:0]   p0_cmd_bl,
  input   [29:0]  p0_cmd_byte_addr,
  output          p0_cmd_empty,
  output          p0_cmd_full,
  input           p0_wr_clk,
  input           p0_wr_en,
  input   [3:0]   p0_wr_mask,
  input   [31:0]  p0_wr_data,
  output          p0_wr_full,
  output          p0_wr_empty,
  output  [6:0]   p0_wr_count,
  output          p0_wr_underrun,
  output          p0_wr_error,
  input           p0_rd_clk,
  input           p0_rd_en,
  output  [31:0]  p0_rd_data,
  output          p0_rd_full,
  output          p0_rd_empty,
  output  [6:0]   p0_rd_count,
  output          p0_rd_overflow,
  output          p0_rd_error,

  input           p1_cmd_clk,
  input           p1_cmd_en,
  input   [2:0]   p1_cmd_instr,
  input   [5:0]   p1_cmd_bl,
  input   [29:0]  p1_cmd_byte_addr,
  output          p1_cmd_empty,
  output          p1_cmd_full,
  input           p1_wr_clk,
  input           p1_wr_en,
  input   [3:0]   p1_wr_mask,
  input   [31:0]  p1_wr_data,
  output          p1_wr_full,
  output          p1_wr_empty,
  output  [6:0]   p1_wr_count,
  output          p1_wr_underrun,
  output          p1_wr_error,
  input           p1_rd_clk,
  input           p1_rd_en,
  output  [31:0]  p1_rd_data,
  output          p1_rd_full,
  output          p1_rd_empty,
  output  [6:0]   p1_rd_count,
  output          p1_rd_overflow,
  output          p1_rd_error,

  input           p2_cmd_clk,
  input           p2_cmd_en,
  input  [2:0]    p2_cmd_instr,
  input  [5:0]    p2_cmd_bl,
  input  [29:0]   p2_cmd_byte_addr,
  output          p2_cmd_empty,
  output          p2_cmd_full,
  input           p2_wr_clk,
  input           p2_wr_en,
  input  [3:0]    p2_wr_mask,
  input  [31:0]   p2_wr_data,
  output          p2_wr_full,
  output          p2_wr_empty,
  output [6:0]    p2_wr_count,
  output          p2_wr_underrun,
  output          p2_wr_error,

  input           p3_cmd_clk,
  input           p3_cmd_en,
  input  [2:0]    p3_cmd_instr,
  input  [5:0]    p3_cmd_bl,
  input  [29:0]   p3_cmd_byte_addr,
  output          p3_cmd_empty,
  output          p3_cmd_full,
  input           p3_wr_clk,
  input           p3_wr_en,
  input  [3:0]    p3_wr_mask,
  input  [31:0]   p3_wr_data,
  output          p3_wr_full,
  output          p3_wr_empty,
  output [6:0]    p3_wr_count,
  output          p3_wr_underrun,
  output          p3_wr_error,

  input           p4_cmd_clk,
  input           p4_cmd_en,
  input  [2:0]    p4_cmd_instr,
  input  [5:0]    p4_cmd_bl,
  input  [29:0]   p4_cmd_byte_addr,
  output          p4_cmd_empty,
  output          p4_cmd_full,
  input           p4_rd_clk,
  input           p4_rd_en,
  output [31:0]   p4_rd_data,
  output          p4_rd_full,
  output          p4_rd_empty,
  output [6:0]    p4_rd_count,
  output          p4_rd_overflow,
  output          p4_rd_error,

  input           p5_cmd_clk,
  input           p5_cmd_en,
  input  [2:0]    p5_cmd_instr,
  input  [5:0]    p5_cmd_bl,
  input  [29:0]   p5_cmd_byte_addr,
  output          p5_cmd_empty,
  output          p5_cmd_full,
  input           p5_rd_clk,
  input           p5_rd_en,
  output [31:0]   p5_rd_data,
  output          p5_rd_full,
  output          p5_rd_empty,
  output [6:0]    p5_rd_count,
  output          p5_rd_overflow,
  output          p5_rd_error


);

artemis_ddr3_base ddr3_base(
  .c3_sys_clk             (clk_333mhz            ),
  .c3_sys_rst_i           (board_rst             ),

  .c3_calib_done          (calibration_done      ),

  .c3_clk0                (usr_clk               ),
  .c3_rst0                (rst                   ),

  .mcb3_dram_dq           (ddr3_dram_dq          ),
  .mcb3_dram_a            (ddr3_dram_a           ),
  .mcb3_dram_ba           (ddr3_dram_ba          ),
  .mcb3_dram_ras_n        (ddr3_dram_ras_n       ),
  .mcb3_dram_cas_n        (ddr3_dram_cas_n       ),
  .mcb3_dram_we_n         (ddr3_dram_we_n        ),
  .mcb3_dram_odt          (ddr3_dram_odt         ),
  .mcb3_dram_reset_n      (ddr3_dram_reset_n     ),
  .mcb3_dram_cke          (ddr3_dram_cke         ),
  .mcb3_dram_dm           (ddr3_dram_dm          ),
  .mcb3_rzq               (ddr3_rzq              ),
  .mcb3_zio               (ddr3_zio              ),
  .mcb3_dram_dqs          (ddr3_dram_dqs         ),
  .mcb3_dram_dqs_n        (ddr3_dram_dqs_n       ),
  .mcb3_dram_ck           (ddr3_dram_ck          ),
  .mcb3_dram_ck_n         (ddr3_dram_ck_n        ),

  .c3_p0_cmd_clk          (p0_cmd_clk            ),
  .c3_p0_cmd_en           (p0_cmd_en             ),
  .c3_p0_cmd_instr        (p0_cmd_instr          ),
  .c3_p0_cmd_bl           (p0_cmd_bl             ),
  .c3_p0_cmd_byte_addr    (p0_cmd_byte_addr      ),
  .c3_p0_cmd_empty        (p0_cmd_empty          ),
  .c3_p0_cmd_full         (p0_cmd_full           ),
  .c3_p0_wr_clk           (p0_wr_clk             ),
  .c3_p0_wr_en            (p0_wr_en              ),
  .c3_p0_wr_mask          (p0_wr_mask            ),
  .c3_p0_wr_data          (p0_wr_data            ),
  .c3_p0_wr_full          (p0_wr_full            ),
  .c3_p0_wr_empty         (p0_wr_empty           ),
  .c3_p0_wr_count         (p0_wr_count           ),
  .c3_p0_wr_underrun      (p0_wr_underrun        ),
  .c3_p0_wr_error         (p0_wr_error           ),
  .c3_p0_rd_clk           (p0_rd_clk             ),
  .c3_p0_rd_en            (p0_rd_en              ),
  .c3_p0_rd_data          (p0_rd_data            ),
  .c3_p0_rd_full          (p0_rd_full            ),
  .c3_p0_rd_empty         (p0_rd_empty           ),
  .c3_p0_rd_count         (p0_rd_count           ),
  .c3_p0_rd_overflow      (p0_rd_overflow        ),
  .c3_p0_rd_error         (p0_rd_error           ),

  .c3_p1_cmd_clk          (p1_cmd_clk            ),
  .c3_p1_cmd_en           (p1_cmd_en             ),
  .c3_p1_cmd_instr        (p1_cmd_instr          ),
  .c3_p1_cmd_bl           (p1_cmd_bl             ),
  .c3_p1_cmd_byte_addr    (p1_cmd_byte_addr      ),
  .c3_p1_cmd_empty        (p1_cmd_empty          ),
  .c3_p1_cmd_full         (p1_cmd_full           ),
  .c3_p1_wr_clk           (p1_wr_clk             ),
  .c3_p1_wr_en            (p1_wr_en              ),
  .c3_p1_wr_mask          (p1_wr_mask            ),
  .c3_p1_wr_data          (p1_wr_data            ),
  .c3_p1_wr_full          (p1_wr_full            ),
  .c3_p1_wr_empty         (p1_wr_empty           ),
  .c3_p1_wr_count         (p1_wr_count           ),
  .c3_p1_wr_underrun      (p1_wr_underrun        ),
  .c3_p1_wr_error         (p1_wr_error           ),
  .c3_p1_rd_clk           (p1_rd_clk             ),
  .c3_p1_rd_en            (p1_rd_en              ),
  .c3_p1_rd_data          (p1_rd_data            ),
  .c3_p1_rd_full          (p1_rd_full            ),
  .c3_p1_rd_empty         (p1_rd_empty           ),
  .c3_p1_rd_count         (p1_rd_count           ),
  .c3_p1_rd_overflow      (p1_rd_overflow        ),
  .c3_p1_rd_error         (p1_rd_error           ),



  .c3_p2_cmd_clk          (p2_cmd_clk            ),
  .c3_p2_cmd_en           (p2_cmd_en             ),
  .c3_p2_cmd_instr        (p2_cmd_instr          ),
  .c3_p2_cmd_bl           (p2_cmd_bl             ),
  .c3_p2_cmd_byte_addr    (p2_cmd_byte_addr      ),
  .c3_p2_cmd_empty        (p2_cmd_empty          ),
  .c3_p2_cmd_full         (p2_cmd_full           ),
  .c3_p2_wr_clk           (p2_wr_clk             ),
  .c3_p2_wr_en            (p2_wr_en              ),
  .c3_p2_wr_mask          (p2_wr_mask            ),
  .c3_p2_wr_data          (p2_wr_data            ),
  .c3_p2_wr_full          (p2_wr_full            ),
  .c3_p2_wr_empty         (p2_wr_empty           ),
  .c3_p2_wr_count         (p2_wr_count           ),
  .c3_p2_wr_underrun      (p2_wr_underrun        ),
  .c3_p2_wr_error         (p2_wr_error           ),
                                                 
  .c3_p3_cmd_clk          (p3_cmd_clk            ),
  .c3_p3_cmd_en           (p3_cmd_en             ),
  .c3_p3_cmd_instr        (p3_cmd_instr          ),
  .c3_p3_cmd_bl           (p3_cmd_bl             ),
  .c3_p3_cmd_byte_addr    (p3_cmd_byte_addr      ),
  .c3_p3_cmd_empty        (p3_cmd_empty          ),
  .c3_p3_cmd_full         (p3_cmd_full           ),
  .c3_p3_wr_clk           (p3_wr_clk             ),
  .c3_p3_wr_en            (p3_wr_en              ),
  .c3_p3_wr_mask          (p3_wr_mask            ),
  .c3_p3_wr_data          (p3_wr_data            ),
  .c3_p3_wr_full          (p3_wr_full            ),
  .c3_p3_wr_empty         (p3_wr_empty           ),
  .c3_p3_wr_count         (p3_wr_count           ),
  .c3_p3_wr_underrun      (p3_wr_underrun        ),
  .c3_p3_wr_error         (p3_wr_error           ),
                                                 
  .c3_p4_cmd_clk          (p4_cmd_clk            ),
  .c3_p4_cmd_en           (p4_cmd_en             ),
  .c3_p4_cmd_instr        (p4_cmd_instr          ),
  .c3_p4_cmd_bl           (p4_cmd_bl             ),
  .c3_p4_cmd_byte_addr    (p4_cmd_byte_addr      ),
  .c3_p4_cmd_empty        (p4_cmd_empty          ),
  .c3_p4_cmd_full         (p4_cmd_full           ),
  .c3_p4_rd_clk           (p4_rd_clk             ),
  .c3_p4_rd_en            (p4_rd_en              ),
  .c3_p4_rd_data          (p4_rd_data            ),
  .c3_p4_rd_full          (p4_rd_full            ),
  .c3_p4_rd_empty         (p4_rd_empty           ),
  .c3_p4_rd_count         (p4_rd_count           ),
  .c3_p4_rd_overflow      (p4_rd_overflow        ),
  .c3_p4_rd_error         (p4_rd_error           ),
                                                 
  .c3_p5_cmd_clk          (p5_cmd_clk            ),
  .c3_p5_cmd_en           (p5_cmd_en             ),
  .c3_p5_cmd_instr        (p5_cmd_instr          ),
  .c3_p5_cmd_bl           (p5_cmd_bl             ),
  .c3_p5_cmd_byte_addr    (p5_cmd_byte_addr      ),
  .c3_p5_cmd_empty        (p5_cmd_empty          ),
  .c3_p5_cmd_full         (p5_cmd_full           ),
  .c3_p5_rd_clk           (p5_rd_clk             ),
  .c3_p5_rd_en            (p5_rd_en              ),
  .c3_p5_rd_data          (p5_rd_data            ),
  .c3_p5_rd_full          (p5_rd_full            ),
  .c3_p5_rd_empty         (p5_rd_empty           ),
  .c3_p5_rd_count         (p5_rd_count           ),
  .c3_p5_rd_overflow      (p5_rd_overflow        ),
  .c3_p5_rd_error         (p5_rd_error           )

);


endmodule
