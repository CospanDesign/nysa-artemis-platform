

module artemis_ddr3 (
  input           clk_333mhz,
  input           board_rst,
  output          calibration_done,
  output          usr_clk,
  output          rst,

  //Memory Interface
  inout  [7:0]    ddr3_dram_dq,
  output [13:0]   ddr3_dram_a,
  output [2:0]    ddr3_dram_ba,
  output          ddr3_dram_ras_n,
  output          ddr3_dram_cas_n,
  output          ddr3_dram_we_n,
  output          ddr3_dram_odt,
  output          ddr3_dram_reset_n,
  output          ddr3_dram_cke,
  output          ddr3_dram_dm,
  inout           ddr3_rzq,
  inout           ddr3_zio,
  inout           ddr3_dram_dqs,
  inout           ddr3_dram_dqs_n,
  output          ddr3_dram_ck,
  output          ddr3_dram_ck_n,

  //Port Interfaces
  input           p0_cmd_clk,
  input           p0_cmd_en,
  input   [2:0]   p0_cmd_instr,
  input   [5:0]   p0_cmd_bl,
  input   [29:0]  p0_cmd_byte_addr,
  output          p0_cmd_empty,
  output          p0_cmd_full,
  input           p0_wr_clk,
  input           p0_wr_en,
  input   [3:0]   p0_wr_mask,
  input   [31:0]  p0_wr_data,
  output          p0_wr_full,
  output          p0_wr_empty,
  output  [6:0]   p0_wr_count,
  output          p0_wr_underrun,
  output          p0_wr_error,
  input           p0_rd_clk,
  input           p0_rd_en,
  output  [31:0]  p0_rd_data,
  output          p0_rd_full,
  output          p0_rd_empty,
  output  [6:0]   p0_rd_count,
  output          p0_rd_overflow,
  output          p0_rd_error,

  input           p1_cmd_clk,
  input           p1_cmd_en,
  input   [2:0]   p1_cmd_instr,
  input   [5:0]   p1_cmd_bl,
  input   [29:0]  p1_cmd_byte_addr,
  output          p1_cmd_empty,
  output          p1_cmd_full,
  input           p1_wr_clk,
  input           p1_wr_en,
  input   [3:0]   p1_wr_mask,
  input   [31:0]  p1_wr_data,
  output          p1_wr_full,
  output          p1_wr_empty,
  output  [6:0]   p1_wr_count,
  output          p1_wr_underrun,
  output          p1_wr_error,
  input           p1_rd_clk,
  input           p1_rd_en,
  output  [31:0]  p1_rd_data,
  output          p1_rd_full,
  output          p1_rd_empty,
  output  [6:0]   p1_rd_count,
  output          p1_rd_overflow,
  output          p1_rd_error,

  input           p2_cmd_clk,
  input           p2_cmd_en,
  input  [2:0]    p2_cmd_instr,
  input  [5:0]    p2_cmd_bl,
  input  [29:0]   p2_cmd_byte_addr,
  output          p2_cmd_empty,
  output          p2_cmd_full,
  input           p2_wr_clk,
  input           p2_wr_en,
  input  [3:0]    p2_wr_mask,
  input  [31:0]   p2_wr_data,
  output          p2_wr_full,
  output          p2_wr_empty,
  output [6:0]    p2_wr_count,
  output          p2_wr_underrun,
  output          p2_wr_error,

  input           p3_cmd_clk,
  input           p3_cmd_en,
  input  [2:0]    p3_cmd_instr,
  input  [5:0]    p3_cmd_bl,
  input  [29:0]   p3_cmd_byte_addr,
  output          p3_cmd_empty,
  output          p3_cmd_full,
  input           p3_wr_clk,
  input           p3_wr_en,
  input  [3:0]    p3_wr_mask,
  input  [31:0]   p3_wr_data,
  output          p3_wr_full,
  output          p3_wr_empty,
  output [6:0]    p3_wr_count,
  output          p3_wr_underrun,
  output          p3_wr_error,

  input           p4_cmd_clk,
  input           p4_cmd_en,
  input  [2:0]    p4_cmd_instr,
  input  [5:0]    p4_cmd_bl,
  input  [29:0]   p4_cmd_byte_addr,
  output          p4_cmd_empty,
  output          p4_cmd_full,
  input           p4_rd_clk,
  input           p4_rd_en,
  output [31:0]   p4_rd_data,
  output          p4_rd_full,
  output          p4_rd_empty,
  output [6:0]    p4_rd_count,
  output          p4_rd_overflow,
  output          p4_rd_error,

  input           p5_cmd_clk,
  input           p5_cmd_en,
  input  [2:0]    p5_cmd_instr,
  input  [5:0]    p5_cmd_bl,
  input  [29:0]   p5_cmd_byte_addr,
  output          p5_cmd_empty,
  output          p5_cmd_full,
  input           p5_rd_clk,
  input           p5_rd_en,
  output [31:0]   p5_rd_data,
  output          p5_rd_full,
  output          p5_rd_empty,
  output [6:0]    p5_rd_count,
  output          p5_rd_overflow,
  output          p5_rd_error


);
endmodule
